module branch_unit #(
    parameter
        WIDTH = 32
) (
    input   [WIDTH-1:0] data_in_1, data_in_2,

    output  reg         branch_en
);
    
endmodule