module RV32I_top_level #(
    parameter
        WIDTH = 32
) (
    input   [WIDTH-1:0] data_in,
    output  [WIDTH-1:0] data_out
);

    wire [WIDTH-1:0]    inst_data;
    
endmodule