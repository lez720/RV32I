module RV32I_top_level #()();