module RV32I_TB;

reg 




endmodule

